netcdf synoptic  {				// synoptic netCDF definition

dimensions:
	recNum = UNLIMITED ;
	rep_type_len = 4;
	stnName_len = 6;
	cloud_levels = 3;
	r_len = 256;

variables:

	char rep_type( recNum, rep_type_len ) ;
		rep_type:long_name = "Report type";
		rep_type:reference = "WMO #306, FM 12-X";
	int wmoId( recNum ) ;
		wmoId:long_name = "WMO Identification number";
		wmoId:_FillValue = -99999;
		wmoId:reference = "systns_upc.tbl Table";
	char stnName( recNum, stnName_len ) ;
		stnName:long_name = "Station Name";
	int time_obs( recNum ) ;
		time_obs:long_name = "time of Observation";
		time_obs:_FillValue = -99999;
		time_obs:units = "seconds since 1970-01-01 00 UTC";
	int time_nominal( recNum ) ;
		time_nominal:long_name = "time nominal";
		time_nominal:_FillValue = -99999;
		time_nominal:units = "seconds since 1970-01-01 00 UTC";
	float Lat( recNum ) ;
		Lat:long_name = "Station latitude";
		Lat:_FillValue = -99999.f;
		Lat:valid_range = -90.0, 90.0;
		Lat:units = "degrees_north";
	float Lon( recNum ) ;
		Lon:long_name = "Station longitude";
		Lon:_FillValue = -99999.f;
		Lon:valid_range = -180.0, 180.0;
		Lon:units = "degrees_east";
	int elev( recNum ) ;
		elev:long_name = "Elevation of station";
		elev:_FillValue = -99999;
		elev:units = "meters";
	int stnType( recNum ) ;
		stnType:long_name = "Type of station operation";
		stnType:_FillValue = -99999;
		stnType:reference = "Table 1860";
	int meanWind( recNum ) ;
		meanWind:long_name = "Highest mean wind speed";
		meanWind:_FillValue = -99999;
		meanWind:reference = "Table 3778";
	int VIS( recNum ) ;
		VIS:long_name = "Horizontal visibility";
		VIS:_FillValue = -99999;
		VIS:reference = "Table 4377";
	int DIR( recNum ) ;
		DIR:long_name = "Wind Direction";
		DIR:_FillValue = -99999;
		DIR:valid_range = 0, 360;
		DIR:units = "degree_true";
	float SPD( recNum ) ;
		SPD:long_name = "Wind Speed";
		SPD:_FillValue = -99999.f;
		SPD:units = "meters/sec";
	float T( recNum ) ;
		T:long_name = "Air Temperature to tenths";
		T:_FillValue = -99999.f;
		T:units = "Celsius";
	int humidity( recNum ) ;
		humidity:long_name = "Humidity";
		humidity:_FillValue = -99999;
		humidity:units = "percent";
	float TD( recNum ) ;
		TD:long_name = "Dew-point Air temperature to tenths";
		TD:_FillValue = -99999.f;
		TD:units = "Celsius";
	float PRES( recNum ) ;
		PRES:long_name = "Station level pressure";
		PRES:_FillValue = -99999.f;
		PRES:units = "hectopascals";
	float SLP( recNum ) ;
		SLP:long_name = "Sea level pressure";
		SLP:_FillValue = -99999.f;
		SLP:units = "hectopascals";
	int char_Ptend( recNum ) ;
		char_Ptend:long_name = "Character Pressure tendency";
		char_Ptend:_FillValue = -99999;
		char_Ptend:reference = "0|1|2|3|4|5|6|7|8 Table 12-5";
		char_Ptend:valid_range = 0, 8;
		char_Ptend:units = "" ;       // dimensionless
	float Ptend( recNum ) ;
		Ptend:long_name = "Change in Pressure in past 3 hours";
		Ptend:_FillValue = -99999.f;
		Ptend:units = "hectopascals";
	float PRECIP_amt( recNum ) ;
		PRECIP_amt:long_name = "Precipitation amount";
		PRECIP_amt:_FillValue = -99999.f;
		PRECIP_amt:units = ".01 meter";
		PRECIP_amt:reference = "Table 3590";
	int PRECIP_period( recNum ) ;
		PRECIP_period:long_name = "Precipitation Period";
		PRECIP_period:_FillValue = -99999;
		PRECIP_period:units = "hours";
		PRECIP_period:reference = "Table 4019";
	int WXpresent( recNum ) ;
		WXpresent:long_name = "Present weather";
		WXpresent:_FillValue = -99999;
		WXpresent:reference = "Manned stn Table 4677, auto Table 4680";
	int WXpast( recNum ) ;
		WXpast:long_name = "Past weather";
		WXpast:_FillValue = -99999;
		WXpast:reference = "Manned stn Table 4561, auto Table 4531";
	int cloudCover( recNum ) ;
		cloudCover:long_name = "Total cloud cover in oktas";
		cloudCover:_FillValue = -99999;
		cloudCover:reference = "Table 2700";
	int cloudLow( recNum ) ;
		cloudLow:long_name = "Lower level clouds";
		cloudLow:_FillValue = -99999;
		cloudLow:reference = "Table 0513";
	int cloudMiddle( recNum ) ;
		cloudMiddle:long_name = "Middle level clouds";
		cloudMiddle:_FillValue = -99999;
		cloudMiddle:reference = "Table 0515";
	int cloudHigh( recNum ) ;
		cloudHigh:long_name = "Higher level clouds";
		cloudHigh:_FillValue = -99999;
		cloudHigh:reference = "Table 0509";
	//int shipTrueDIR( recNum ) ;
		//shipTrueDIR:long_name = "Ship's True direction";
		//shipTrueDIR:_FillValue = -99999;
		//shipTrueDIR:reference = "Table 0700";
	//int shipAvgSPD( recNum ) ;
		//shipAvgSPD:long_name = "Ship's Avg speed";
		//shipAvgSPD:_FillValue = -99999;
		//shipAvgSPD:reference = "Table 4451";
	float Tw( recNum ) ;
		Tw:long_name = "Water Temperature to tenths";
		Tw:_FillValue = -99999.f;
		Tw:units = "Celsius";
	int Pwa( recNum ) ;
		Pwa:long_name = "Period of waves";
		Pwa:_FillValue = -99999;
		Pwa:units = "seconds";
	int Hwa( recNum ) ;
		Hwa:long_name = "Height of waves";
		Hwa:_FillValue = -99999;
		Hwa:units = "meters";
	float Hwa_tenths( recNum ) ;
		Hwa_tenths:long_name = "Height of waves";
		Hwa_tenths:_FillValue = -99999.f;
		Hwa_tenths:units = "meters";
	int swellDIR1( recNum ) ;
		swellDIR1:long_name = "Direction of swells";
		swellDIR1:_FillValue = -99999;
		swellDIR1:units = "degrees";
	float Ps1( recNum ) ;
		Ps1:long_name = "Period of swells";
		Ps1:_FillValue = -99999.f;
		Ps1:units = "seconds";
	float Hs1( recNum ) ;
		Hs1:long_name = "Height of swells";
		Hs1:_FillValue = -99999.f;
		Hs1:units = "meters";
	//int swellDIR2( recNum ) ;
		//swellDIR2:long_name = "Direction of swells";
		//swellDIR2:_FillValue = -99999;
		//swellDIR2:units = "degree_true";
	//float Ps2( recNum ) ;
		//Ps2:long_name = "Period of swells";
		//Ps2:_FillValue = -99999.f;
		//Ps2:units = "seconds";
	//float Hs2( recNum ) ;
		//Hs2:long_name = "Height of swells";
		//Hs2:_FillValue = -99999.f;
		//Hs2:units = "meters";
	//int iceType( recNum ) ;
		//iceType:long_name = "Type of Ice build up";
		//iceType:_FillValue = -99999;
		//iceType:reference = "Table 1751";
	//int iceThick( recNum ) ;
		//iceThick:long_name = "Ice thickness";
		//iceThick:_FillValue = -99999;
		//iceThick:units = "centimeters";
	//int iceRate( recNum ) ;
		//iceRate:long_name = "Rate of Ice build up";
		//iceRate:_FillValue = -99999;
		//iceRate:reference = "Table 3551";
	float Tb( recNum ) ;
		Tb:long_name = "Web Bulb Temperature";
		Tb:_FillValue = -99999.f;
		Tb:units = "Celsius";
	int ICE( recNum ) ;
		ICE:long_name = "Sea ice or ice of land origin";
		ICE:_FillValue = -99999;
	//int iceConcen( recNum ) ;
		//iceConcen:long_name = "Ice concentration";
		//iceConcen:_FillValue = -99999;
		//iceConcen:reference = "Table 0639";
	//int iceStage( recNum ) ;
		//iceStage:long_name = "Stage of development";
		//iceStage:_FillValue = -99999;
		//iceStage:reference = "Table 3739";
	//int iceLand( recNum ) ;
		//iceLand:long_name = "Ice of Land origin";
		//iceLand:_FillValue = -99999;
		//iceLand:reference = "Table 0439";
	//int iceEdge( recNum ) ;
		//iceEdge:long_name = "True bearing of Ice Edge";
		//iceEdge:_FillValue = -99999;
		//iceEdge:reference = "Table 0739";
	//int iceSituation( recNum ) ;
		//iceSituation:long_name = "Present Ice Situation";
		//iceSituation:_FillValue = -99999;
		//iceSituation:reference = "Table 5239";
	float Tmax( recNum ) ;
		Tmax:long_name = "Max Air Temperature to tenths";
		Tmax:_FillValue = -99999.f;
		Tmax:units = "Celsius";
	float Tmin( recNum ) ;
		Tmin:long_name = "Min Air Temperature to tenths";
		Tmin:_FillValue = -99999.f;
		Tmin:units = "Celsius";
	int groundState( recNum ) ;
		groundState:long_name = "State of ground";
		groundState:_FillValue = -99999;
		groundState:reference = "Table 0975";
	int snowDepth( recNum ) ;
		snowDepth:long_name = "Snow depth";
		snowDepth:_FillValue = -99999;
		snowDepth:units = "centimeters";
		snowDepth:reference = "Table 3889";
	float PRECIP_amt24( recNum ) ;
		PRECIP_amt24:long_name = "Precipitation amount last 24 hours";
		PRECIP_amt24:_FillValue = -99999.f;
		PRECIP_amt24:units = ".01 meter";
	int cloudObsured( recNum, cloud_levels ) ;
		cloudObsured:long_name = "Total cloud cover in oktas";
		cloudObsured:_FillValue = -99999;
		cloudObsured:reference = "Table 2700";
	int cloudGenus( recNum, cloud_levels ) ;
		cloudGenus:long_name = "Cloud genus";
		cloudGenus:_FillValue = -99999;
		cloudGenus:reference = "Table 0500";
	int cloudHeight( recNum, cloud_levels ) ;
		cloudHeight:long_name = "Cloud Height in meters";
		cloudHeight:_FillValue = -99999;
		cloudHeight:reference = "Table 1677";
	char report( recNum, r_len ) ;
		report:long_name = "Originial report";
		report:reference = "max length 256";

	:title = "SYNOPTIC definition";
	:version = 1.1;

//	In general:
//	
//	The syn2nc decoder is dependant on the netCDF variables names 
//	because it reads the cdl file to determine the variables to be
//	included in the netcdf file.  A user can comment out or delete
//	variables not to be included in the output file with exceptions,
//	the variables 'rep_type', 'wmoId' must be included.
//	The WMO Manual on Codes #306 FM 12-X and FM 18-IX was used for some 
//	variable definitions and all tables references are also from the same 
//	manual.
//	
//	Units must be compatible with UDUNITS and consistent for a given 
//	variable (ie. all temperatures written out in degrees C, even though
//	they are reported in C or F). That's why the "units" attribute is
//	critical for numeric variables that may be used in calculations.
//	
} 
